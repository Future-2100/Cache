
package core_pkg;

`include "core_trans.sv"

`include "core_generator.sv"

`include "core_driver.sv"

`include "core_monitor.sv"

`include "core_agent.sv"

endpackage

