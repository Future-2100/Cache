
package cache_pkg;

import core_pkg::*;

import  axi_pkg::*;

import  rpt_pkg::*;

`include "cache_checker.sv"

`include "cache_coverage.sv"

`include "cache_env.sv"

`include "base_test.sv"

endpackage:cache_pkg

