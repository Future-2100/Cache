
package axi_pkg;

`include "axi_trans.sv"

`include "axi_driver.sv"

`include "axi_generator.sv"

endpackage
